// TargetMatrixBitMap File 
// A two level bitmap. dosplaying Target on the screen FWbruary  2021  
// (c) Technion IIT, Department of Electrical Engineering 2021 



module	TargetMatrixBitMap	(	
					input	logic	clk,
					input	logic	resetN,
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY,
					input	logic	InsideRectangle, //input that the pixel is within a bracket 

					output	logic	drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[7:0] RGBout  //rgb value from the bitmap 
 ) ;
 

// Size represented as Number of X and Y bits 
localparam logic [7:0] TRANSPARENT_ENCODING = 8'h00 ;// RGB value in the bitmap representing a transparent pixel 
 /*  end generated by the tool */


// the screen is 640*480  or  10 * 15 squares of 32*32  bits ,  we wiil round up to 16*16 and use only the top left 10*15 pixels  
// this is the bitmap  of the maze , if there is a one  the na whole 32*32 rectange will be drawn on the screen 
// all numbers here are hard coded to simplify the  understanding 


logic [0:7] [0:7]  MazeBiMapMask= 
{8'b	00000000,
8'b	00000000,
8'b	00000000,
8'b	00000000,
8'b	00000000,
8'b	00000000,
8'b	10000000
};
 
 logic[0:63][0:63][7:0] object_colors = {
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h00,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h01,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h01,8'h01,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h42,8'h01,8'h01,8'h00,8'h00},
	{8'h00,8'h01,8'h01,8'h42,8'h42,8'h8b,8'h8b,8'h8b,8'h8a,8'h8a,8'h8a,8'h8a,8'h8b,8'h8b,8'h8b,8'h8b,8'h8a,8'h8a,8'h8a,8'h8a,8'h8a,8'h8a,8'h8a,8'h8b,8'h8b,8'h8b,8'h8a,8'h8b,8'h8b,8'h8b,8'h8b,8'h8b,8'h8b,8'h8b,8'h8b,8'h8a,8'h8b,8'h8b,8'h8b,8'h8b,8'h8b,8'h8a,8'h8a,8'h8b,8'h8b,8'h8a,8'h8b,8'h8b,8'h8b,8'h8b,8'h8b,8'h8b,8'h8b,8'h8b,8'h8b,8'h8a,8'h8b,8'h8b,8'h8b,8'h42,8'h42,8'h01,8'h00,8'h00},
	{8'h01,8'h01,8'h42,8'h42,8'h8b,8'hd3,8'h93,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'h8b,8'h42,8'h42,8'h01,8'h00},
	{8'h01,8'h42,8'h42,8'h42,8'h42,8'h01,8'h01,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'h49,8'hd3,8'h41,8'h00,8'h00,8'h00,8'h40,8'h40,8'h89,8'h89,8'h89,8'h89,8'h89,8'h89,8'h89,8'h89,8'h89,8'h40,8'h00,8'h00,8'h00,8'h00,8'h00,8'h49,8'hd3,8'h41,8'h40,8'h41,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'h89,8'h00,8'h00,8'h00,8'h00,8'h01,8'h01,8'h42,8'h42,8'h42,8'h42,8'h01},
	{8'h42,8'h43,8'h43,8'h8b,8'h42,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h41,8'hd3,8'h41,8'h00,8'h00,8'h00,8'h40,8'h40,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h40,8'h00,8'h00,8'h00,8'h00,8'h00,8'h49,8'hd3,8'h41,8'h40,8'h89,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd1,8'h89,8'h89,8'h8a,8'h8a,8'h49,8'h01,8'h8a,8'h8b,8'h42,8'h42,8'h42},
	{8'h42,8'h42,8'h42,8'hd3,8'h8a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h49,8'hdb,8'h40,8'h00,8'h00,8'h00,8'h40,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h40,8'h00,8'h00,8'h00,8'h00,8'h49,8'hd3,8'h40,8'h89,8'hd2,8'hd2,8'hd1,8'hd1,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hdb,8'hdb,8'h92,8'h00,8'h8a,8'h8b,8'h42,8'h42,8'h42},
	{8'h8b,8'h8a,8'h01,8'h41,8'h4a,8'h8a,8'h00,8'h00,8'h00,8'h00,8'h89,8'h91,8'h91,8'h91,8'h91,8'h49,8'h00,8'h00,8'h00,8'h41,8'hd3,8'h40,8'h00,8'h00,8'h40,8'h88,8'h89,8'hd1,8'hd1,8'hc8,8'h88,8'h88,8'h88,8'hd1,8'hd1,8'hd1,8'h88,8'h40,8'h40,8'h00,8'h00,8'h00,8'h49,8'hdb,8'h92,8'hd2,8'hd2,8'hd1,8'hd1,8'hd1,8'hd2,8'hd2,8'hd1,8'hd2,8'hd2,8'hd2,8'hd3,8'hd3,8'h92,8'h49,8'h41,8'h01,8'h8b,8'h8b},
	{8'h8b,8'h8b,8'h00,8'h00,8'h41,8'h89,8'h49,8'h49,8'h49,8'h49,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'h91,8'h48,8'h00,8'h00,8'h41,8'hd3,8'h40,8'h00,8'h40,8'h88,8'h89,8'hd1,8'hd2,8'hd2,8'hd1,8'hc8,8'h88,8'hd1,8'hd1,8'hd2,8'hd1,8'hd1,8'h88,8'h40,8'h40,8'h00,8'h00,8'h49,8'hdb,8'h8a,8'hd1,8'hd1,8'hc8,8'hd1,8'hd1,8'hd2,8'hd1,8'hd1,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'h8a,8'h40,8'h00,8'h00,8'hd3,8'h8b},
	{8'h8b,8'h8b,8'h00,8'h00,8'h00,8'h00,8'hd2,8'hdb,8'hd2,8'hd2,8'hd2,8'hd2,8'hd1,8'hc9,8'hd1,8'hd2,8'hd2,8'h40,8'h00,8'h41,8'hdb,8'h49,8'h40,8'h88,8'h88,8'hd1,8'hd2,8'hda,8'hd2,8'hda,8'hd1,8'h88,8'hda,8'hd2,8'hd2,8'hd2,8'hd2,8'hc9,8'h88,8'h88,8'h40,8'h00,8'h49,8'hd3,8'h40,8'h80,8'hc9,8'hc8,8'hc9,8'hc9,8'hd1,8'hc9,8'hd1,8'hd2,8'hd2,8'hd2,8'hd2,8'hca,8'h40,8'h00,8'h00,8'h00,8'hd3,8'h8b},
	{8'h8b,8'h8b,8'h00,8'h00,8'h00,8'h40,8'hd2,8'hda,8'hd2,8'hd2,8'hd2,8'hd2,8'hd1,8'hd1,8'hd1,8'hd1,8'hd2,8'h89,8'h40,8'h41,8'hdb,8'h89,8'h88,8'h88,8'hc9,8'hd1,8'hda,8'hda,8'hda,8'hda,8'hd2,8'h91,8'hdb,8'hda,8'hda,8'hd2,8'hd2,8'hd1,8'h88,8'h88,8'h89,8'h40,8'h49,8'hd3,8'h40,8'h88,8'hd1,8'hc8,8'hc8,8'hc8,8'hc9,8'hc8,8'hc9,8'hc9,8'hc9,8'hc9,8'hc9,8'hc9,8'h80,8'h40,8'h40,8'h40,8'hd3,8'h8b},
	{8'h8b,8'h8b,8'h00,8'h00,8'h00,8'h48,8'hd2,8'hd2,8'hd2,8'hd1,8'hd1,8'hd2,8'hd1,8'hd1,8'hd1,8'hd1,8'hd2,8'h92,8'h40,8'h41,8'hda,8'hd2,8'hd1,8'h88,8'hd1,8'hd2,8'hd2,8'hda,8'hdb,8'hdb,8'hd2,8'hda,8'hd2,8'hdb,8'hda,8'hd2,8'hd2,8'hd1,8'hd1,8'h88,8'hd2,8'h89,8'h89,8'hd3,8'h40,8'h48,8'hc9,8'h80,8'h80,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc1,8'h80,8'h40,8'h40,8'hd3,8'h8b},
	{8'h8b,8'h8a,8'h00,8'h00,8'h89,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd1,8'hd1,8'hd1,8'hc9,8'hc8,8'hc9,8'h89,8'h40,8'h00,8'h49,8'hda,8'hd2,8'hd1,8'h88,8'h88,8'hd1,8'hd2,8'hda,8'hdb,8'h89,8'h40,8'hd2,8'h00,8'hdb,8'hda,8'hd2,8'hd2,8'hc9,8'h88,8'h88,8'hd2,8'hd2,8'hd2,8'hd2,8'h40,8'h00,8'h40,8'h80,8'hc9,8'hc9,8'hc0,8'hc9,8'hc9,8'hc0,8'hc0,8'hc9,8'hc9,8'hc0,8'hd2,8'hc9,8'h40,8'h40,8'hd3,8'h8b},
	{8'h8b,8'hcb,8'h40,8'h40,8'h80,8'hc9,8'hd1,8'hc9,8'hc9,8'hc9,8'hc9,8'hc9,8'hc9,8'hc8,8'hc8,8'hc9,8'h89,8'h40,8'h00,8'h49,8'hda,8'hd2,8'hd1,8'h88,8'h88,8'hd1,8'hd2,8'hda,8'hda,8'h89,8'h89,8'hd2,8'h48,8'hda,8'hda,8'hd2,8'hd2,8'h89,8'h88,8'h88,8'hd2,8'hd2,8'hd2,8'hd2,8'h48,8'h40,8'h40,8'h80,8'hc9,8'hc9,8'hc0,8'hc9,8'hc8,8'hc0,8'hc0,8'hc9,8'hc8,8'hc0,8'hc9,8'h89,8'h40,8'h40,8'hd3,8'h8b},
	{8'h8b,8'hd3,8'h81,8'h80,8'h80,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'hc9,8'hd2,8'h00,8'h40,8'h89,8'hd2,8'hd2,8'hd1,8'h88,8'h88,8'hd1,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hda,8'hd2,8'h89,8'h88,8'h88,8'hd2,8'hd2,8'hd2,8'hd2,8'h89,8'h40,8'h40,8'h80,8'h80,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'h80,8'h40,8'h40,8'hd3,8'h8b},
	{8'h8b,8'hcb,8'h81,8'hc9,8'hc9,8'hc0,8'hc9,8'hc0,8'hc0,8'hc0,8'hc9,8'hc9,8'hc0,8'hc9,8'hc0,8'h80,8'h40,8'h00,8'h40,8'h89,8'hd2,8'hd2,8'hd2,8'hd1,8'hd1,8'hd2,8'hd2,8'hd2,8'hd2,8'hd1,8'h88,8'h88,8'hc9,8'hd2,8'hd2,8'hd2,8'hd2,8'hd1,8'hd1,8'hd1,8'hd2,8'hd1,8'hd1,8'hd2,8'h89,8'h40,8'h40,8'h88,8'hc8,8'hc8,8'hc8,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'h40,8'h40,8'h40,8'hd3,8'h8b},
	{8'h8b,8'hcb,8'h81,8'hc9,8'hc0,8'hc0,8'hc9,8'hc0,8'hc0,8'hc0,8'hc9,8'hc0,8'hc0,8'hc9,8'hc0,8'h80,8'h40,8'h40,8'h88,8'h89,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd1,8'hd1,8'hd1,8'hd1,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd1,8'hd1,8'hd2,8'h89,8'h80,8'h80,8'h88,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc0,8'hc8,8'hc8,8'hc0,8'hc8,8'h80,8'h40,8'h00,8'hd3,8'h8b},
	{8'h8b,8'hcb,8'h80,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'h40,8'h48,8'h88,8'h89,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'h89,8'h88,8'h88,8'h88,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'h88,8'h88,8'h40,8'h00,8'hd3,8'h8b},
	{8'h8b,8'hd3,8'h81,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc8,8'hc8,8'hc0,8'h80,8'h40,8'h88,8'h88,8'hc9,8'hd2,8'hd2,8'hd2,8'hd1,8'hd1,8'hc9,8'hc9,8'hc9,8'hd1,8'hc9,8'hc9,8'hc9,8'hc9,8'hc9,8'hc9,8'hd1,8'hc9,8'hd1,8'hd1,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'h89,8'h88,8'h88,8'h88,8'h88,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h40,8'h00,8'hd3,8'h8b},
	{8'h8b,8'hd3,8'h81,8'hc0,8'hc8,8'hc0,8'hc0,8'hc8,8'hc0,8'hc0,8'hc0,8'hc8,8'hc8,8'hc8,8'hc8,8'h80,8'h40,8'h88,8'h88,8'hc9,8'hd2,8'hd2,8'hd2,8'hd1,8'h89,8'hc9,8'h89,8'h89,8'hc9,8'hc9,8'h89,8'h89,8'h89,8'h89,8'h89,8'h89,8'h89,8'h89,8'hd1,8'hd1,8'hd2,8'hd2,8'hd2,8'hd2,8'h89,8'h88,8'h88,8'hc8,8'h88,8'h88,8'hc8,8'hc8,8'hc8,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h40,8'h00,8'hd3,8'h8b},
	{8'h8b,8'hd3,8'h80,8'h88,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'h88,8'h88,8'h88,8'h88,8'h89,8'hda,8'hd2,8'hd1,8'h89,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd1,8'h89,8'hd1,8'hd2,8'hd2,8'hd2,8'h89,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'hc8,8'hc8,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h40,8'h00,8'hd3,8'h8b},
	{8'h8b,8'hd3,8'h89,8'h88,8'h88,8'hc8,8'hc8,8'h88,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'h88,8'h88,8'h88,8'h88,8'h88,8'h89,8'hd2,8'hd1,8'hd1,8'hd1,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd2,8'h89,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h48,8'h40,8'h00,8'hd3,8'h8b},
	{8'h8b,8'hd3,8'h89,8'h88,8'h88,8'h88,8'h88,8'h88,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'hc9,8'hd2,8'h89,8'hc9,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd1,8'h88,8'h88,8'hc9,8'hd2,8'h89,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'hc8,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h40,8'h00,8'h00,8'hd3,8'h8b},
	{8'h8b,8'hd3,8'h89,8'h88,8'hc8,8'hc8,8'h88,8'h88,8'hc8,8'hc8,8'hc8,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'hc9,8'hd2,8'hc9,8'hc9,8'hd1,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd1,8'h88,8'h88,8'hc9,8'hd2,8'h89,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h00,8'h00,8'h00,8'h00,8'hd3,8'h8b},
	{8'h8b,8'hd3,8'h89,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'hc9,8'hd2,8'hc8,8'hc8,8'hc8,8'hd1,8'hd1,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd1,8'hc9,8'hc8,8'h88,8'h88,8'hc9,8'hd2,8'h89,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h48,8'h40,8'h00,8'h00,8'h00,8'h00,8'hd3,8'h8b},
	{8'h8b,8'hd3,8'h89,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'hc9,8'hd1,8'hc8,8'h88,8'h88,8'h88,8'hd1,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hc9,8'h88,8'h88,8'h88,8'h88,8'hc8,8'hd2,8'hc9,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h40,8'h00,8'h00,8'h00,8'h00,8'h00,8'h93,8'h8a},
	{8'h41,8'h41,8'h40,8'h40,8'h40,8'h40,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'hc8,8'hc8,8'h88,8'h88,8'h88,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'h88,8'h88,8'h88,8'h88,8'h88,8'hc8,8'hc9,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h40,8'h40,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h41,8'h41},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h40,8'h40,8'h40,8'h40,8'h40,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'hc8,8'hc8,8'hc8,8'hc8,8'h88,8'hc8,8'hc8,8'h88,8'hc8,8'hc8,8'hc8,8'hc8,8'h88,8'hc8,8'h88,8'h88,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h80,8'h40,8'h40,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h40,8'h40,8'h40,8'h80,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h40,8'h40,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h41,8'h41,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h40,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'hc8,8'hd1,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc9,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h40,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h49,8'h41},
	{8'h8b,8'h8a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h40,8'h88,8'hc8,8'hc8,8'h88,8'h88,8'h88,8'h88,8'h88,8'hc9,8'hd2,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hd2,8'h88,8'h88,8'h88,8'h88,8'h88,8'h40,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h93,8'h8a},
	{8'h8b,8'h8b,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h88,8'h88,8'hc8,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'hc9,8'hd2,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hd1,8'hd2,8'h89,8'h88,8'h88,8'h88,8'hc8,8'h88,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd3,8'h8b},
	{8'h8b,8'h8b,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h40,8'h88,8'hc8,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'hc9,8'hd2,8'hd0,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hd1,8'hd2,8'h89,8'h88,8'h88,8'h88,8'hc8,8'h88,8'h40,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd3,8'h8b},
	{8'h8b,8'h93,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h40,8'hc9,8'hc8,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h89,8'hd2,8'hd0,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hd1,8'hd2,8'h89,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h40,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd3,8'h8b},
	{8'h8b,8'h8b,8'h00,8'h00,8'h00,8'h00,8'h00,8'h40,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'hc9,8'hd2,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hd2,8'h89,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h40,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd3,8'h8b},
	{8'h8b,8'h8b,8'h00,8'h00,8'h00,8'h00,8'h00,8'h88,8'hc8,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'hc9,8'hd2,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hd2,8'h89,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h40,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd3,8'h8b},
	{8'h8b,8'h8b,8'h00,8'h00,8'h00,8'h00,8'h00,8'h88,8'hc8,8'hc8,8'hc8,8'hc8,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'hc9,8'hd2,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hd1,8'hd2,8'h89,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h48,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd3,8'h8b},
	{8'h8b,8'h8b,8'h00,8'h00,8'h00,8'h00,8'h00,8'h88,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'h88,8'hc8,8'hc8,8'h88,8'h88,8'h88,8'hc9,8'hd2,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hd2,8'h89,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'hc8,8'hc8,8'h88,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd3,8'h8b},
	{8'h8b,8'h8b,8'h00,8'h00,8'h00,8'h00,8'h00,8'h88,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'h88,8'h88,8'hc9,8'hd2,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hd2,8'h89,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'hc8,8'h88,8'h40,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd3,8'h8b},
	{8'h8b,8'h93,8'h00,8'h00,8'h00,8'h00,8'h00,8'h88,8'hc8,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc8,8'hc9,8'hd2,8'hc8,8'h88,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'h88,8'hc8,8'hd2,8'h89,8'h88,8'h88,8'h88,8'h88,8'hc8,8'hc8,8'h88,8'h88,8'h88,8'h89,8'h40,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd3,8'h8b},
	{8'h8b,8'h93,8'h00,8'h00,8'h00,8'h00,8'h40,8'h80,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc9,8'hd2,8'hc8,8'h88,8'h88,8'h88,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'h88,8'h88,8'h88,8'hc8,8'hd2,8'h89,8'h88,8'h88,8'h88,8'h88,8'hc8,8'hc8,8'hc8,8'h88,8'h88,8'h89,8'h40,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd3,8'h8b},
	{8'h8b,8'h8b,8'h00,8'h00,8'h00,8'h40,8'h80,8'h80,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'h80,8'hc9,8'hd2,8'hc8,8'h88,8'h88,8'h88,8'h88,8'h88,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'hc8,8'hd2,8'h89,8'h88,8'h88,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc8,8'hc9,8'h40,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd3,8'h8b},
	{8'h8b,8'h8b,8'h00,8'h00,8'h00,8'h40,8'h80,8'hc9,8'hc9,8'hc0,8'hc9,8'hc8,8'hc0,8'hc0,8'hc9,8'hc9,8'hc0,8'hc9,8'hc9,8'hc9,8'hd2,8'h89,8'h40,8'h40,8'h40,8'h40,8'h40,8'h88,8'hc8,8'h88,8'h88,8'hc8,8'h88,8'hc8,8'hc8,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'h88,8'hc9,8'hd2,8'hc9,8'h88,8'hc0,8'hc8,8'hc8,8'hc0,8'hc0,8'hc0,8'hc8,8'hc8,8'hc9,8'h40,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd3,8'h8b},
	{8'h8b,8'h8b,8'h00,8'h00,8'h00,8'h40,8'h80,8'hc9,8'hc9,8'hc0,8'hc9,8'hc0,8'hc0,8'hc0,8'hc9,8'hc1,8'hc0,8'hc9,8'hc1,8'hc9,8'hd2,8'h89,8'h40,8'h00,8'h00,8'h00,8'h00,8'h40,8'h40,8'h40,8'h40,8'h40,8'h40,8'h40,8'h40,8'h40,8'h40,8'h40,8'h40,8'h40,8'h88,8'h88,8'hc9,8'hd2,8'hc9,8'h80,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'h40,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd3,8'h8b},
	{8'h8b,8'h93,8'h00,8'h00,8'h00,8'h40,8'h80,8'h80,8'h80,8'h80,8'hc0,8'hc0,8'h80,8'h80,8'hc0,8'hc0,8'h80,8'h80,8'h80,8'hc9,8'hd2,8'h89,8'h40,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h40,8'h88,8'h88,8'hc9,8'hd2,8'h89,8'h80,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'h80,8'h80,8'h40,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd3,8'h8b},
	{8'h8b,8'h93,8'h00,8'h00,8'h00,8'h40,8'hc9,8'hc9,8'hc9,8'hc9,8'hc9,8'hc9,8'hc9,8'hc9,8'hc9,8'hc9,8'hc9,8'hc9,8'hc9,8'hd2,8'hd2,8'hd2,8'h49,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h40,8'h80,8'hc9,8'hd2,8'hd2,8'hc9,8'hc0,8'hc9,8'hc0,8'hc0,8'hc0,8'hc9,8'hc0,8'hc0,8'hc9,8'h80,8'h40,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd3,8'h8b},
	{8'h8b,8'h8b,8'h00,8'h00,8'h00,8'h89,8'hd2,8'hd2,8'hd2,8'hd2,8'hd1,8'hd2,8'hd2,8'hd1,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd3,8'hd2,8'h89,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h40,8'h89,8'hd2,8'hd2,8'hc9,8'hc0,8'hc9,8'hc0,8'hc0,8'hc0,8'hc9,8'hc0,8'hc0,8'hc9,8'hc0,8'h40,8'h00,8'h41,8'h00,8'h00,8'h00,8'hd3,8'h8b},
	{8'h8b,8'h8b,8'h00,8'h00,8'h49,8'h92,8'hd2,8'hd2,8'hd1,8'hd2,8'hc9,8'hd1,8'hd2,8'h89,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd3,8'hdb,8'hd2,8'h49,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h40,8'h89,8'hd2,8'hc9,8'h81,8'h80,8'hc1,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc9,8'h80,8'h40,8'h00,8'h8a,8'h00,8'h00,8'h00,8'hd3,8'h8b},
	{8'h8b,8'h8b,8'h00,8'h49,8'h49,8'h89,8'h89,8'h49,8'h49,8'h89,8'h48,8'h49,8'h89,8'h40,8'h89,8'h89,8'h89,8'h89,8'h89,8'h92,8'hdb,8'h92,8'h40,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h40,8'h89,8'hd2,8'h89,8'h89,8'hc9,8'hc9,8'hc9,8'hc9,8'hc9,8'hc9,8'hc9,8'hc9,8'hc9,8'hc9,8'h89,8'h49,8'h89,8'h49,8'h41,8'h00,8'hd3,8'h8b},
	{8'h8b,8'h8b,8'h01,8'h92,8'h49,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h49,8'hdb,8'h40,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h41,8'hd3,8'hc9,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'h00,8'h49,8'h8a,8'h41,8'hcb,8'h8b},
	{8'h42,8'h8a,8'hd3,8'h41,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h49,8'hd3,8'h41,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h41,8'hd3,8'hd3,8'hd2,8'hd2,8'hd2,8'hd2,8'hd2,8'h89,8'hd2,8'hd1,8'hc9,8'hd2,8'h8a,8'hd2,8'hd2,8'h00,8'h00,8'h49,8'hd3,8'h8a,8'h42},
	{8'h42,8'h8a,8'hd3,8'h4a,8'h41,8'h41,8'h41,8'h41,8'h41,8'h41,8'h41,8'h41,8'h41,8'h41,8'h41,8'h41,8'h41,8'h41,8'h41,8'h4a,8'hd3,8'h49,8'h41,8'h41,8'h41,8'h41,8'h41,8'h41,8'h41,8'h41,8'h41,8'h41,8'h41,8'h41,8'h41,8'h41,8'h41,8'h41,8'h41,8'h41,8'h41,8'h41,8'h8a,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd2,8'h8a,8'hd3,8'hd2,8'hca,8'hd3,8'hca,8'hd2,8'hd3,8'h41,8'h41,8'h4a,8'hd3,8'h42,8'h42},
	{8'h01,8'h42,8'h42,8'hcb,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'hd3,8'h8b,8'h42,8'h42,8'h01},
	{8'h01,8'h01,8'h42,8'h82,8'h8a,8'h8a,8'h8a,8'h8a,8'h8a,8'h8a,8'h8a,8'h8b,8'h8b,8'h8b,8'h8b,8'h8b,8'h8b,8'h8b,8'h8b,8'h8b,8'h8b,8'h8a,8'h8a,8'h8a,8'h8a,8'h8a,8'h8a,8'h8a,8'h8a,8'h8a,8'h8a,8'h8a,8'h8a,8'h8a,8'h8a,8'h8a,8'h8a,8'h8a,8'h8a,8'h8a,8'h8a,8'h8a,8'h8a,8'h8b,8'h8b,8'h8b,8'h8b,8'h8b,8'h8b,8'h8b,8'h8b,8'h8b,8'h8b,8'h8a,8'h8a,8'h8a,8'h8a,8'h8a,8'h8a,8'h8a,8'h82,8'h42,8'h01,8'h01}};

 
 
//////////--------------------------------------------------------------------------------------------------------------= 
//hit bit map has one bit per edge:  hit_colors[3:0] =   {Left, Top, Right, Bottom}	 
//there is one bit per edge, in the corner two bits are set  
 logic [0:3] [0:3] [3:0] hit_colors = 
		   {16'hC446,     
			16'h8C62,    
			16'h8932, 
			16'h9113}; 
// pipeline (ff) to get the pixel color from the array 	 

//==----------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		RGBout <=	8'h00;
	end
	else begin
		RGBout <= TRANSPARENT_ENCODING ; // default 

		if ((InsideRectangle == 1'b1 )		& 	// only if inside the external bracket 
		   (MazeBiMapMask[offsetY[8:6] ][offsetX[8:6]] == 1'b1 )) // take bits 5,6,7,8,9,10 from address to select  position in the maze    
						RGBout <= object_colors[offsetY[5:0]][offsetX[5:0]] ; 
		end 
end

//==----------------------------------------------------------------------------------------------------------------=
// decide if to draw the pixel or not 
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap   
endmodule