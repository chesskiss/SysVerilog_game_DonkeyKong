// (c) Technion IIT, Department of Electrical Engineering 2021 
//-- Alex Grinshpun Apr 2017
//-- Dudy Nov 13 2017
// SystemVerilog version Alex Grinshpun May 2018
// coding convention dudy December 2018
// updaed Eyal Lev Feb 2021


module	rope_moveCollision	(	
 
					input	logic	clk,
					input	logic	resetN,
					input	logic	startOfFrame,  // short pulse every start of frame 30Hz 
					//input logic singleHit,  //collision if smiley hits an object 
					
					output	 logic  [10:0]	rope_speed,	
					output	 logic signed 	[10:0]	topLeftX, // output the top left corner 
					output	 logic signed	[10:0]	topLeftY  // can be negative , if the object is partliy outside
				  
				 
);


// a module used to generate the  ball trajectory.  

parameter int INITIAL_X = 192;
parameter int INITIAL_Y = 64;//128
parameter int INITIAL_X_SPEED = 20;
parameter int NEGETIVE_X_SPEED = -20;
parameter int INITIAL_Y_SPEED = 0;
parameter int MAX_Y_SPEED = 230;



const int	FIXED_POINT_MULTIPLIER	=	64;
// FIXED_POINT_MULTIPLIER is used to enable working with integers in high resolution so that 
// we do all calculations with topLeftX_FixedPoint to get a resolution of 1/64 pixel in calcuatuions,
// we devide at the end by FIXED_POINT_MULTIPLIER which must be 2^n, to return to the initial proportions
const int	x_FRAME_SIZE	=	575 * FIXED_POINT_MULTIPLIER; // note it must be 2^n //639 ?
//const int	y_FRAME_SIZE	=	479 * FIXED_POINT_MULTIPLIER;
const int	bracketOffset =	30;
const int   OBJECT_WIDTH_X = 32;

int Xspeed, topLeftX_FixedPoint; // local parameters 
int Yspeed, topLeftY_FixedPoint;

assign rope_speed = Xspeed;

//////////--------------------------------------------------------------------------------------------------------------=
//  calculation 0f Y Axis speed using gravity or colision

always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin 
		topLeftY_FixedPoint	<= INITIAL_Y * FIXED_POINT_MULTIPLIER;
	end 
end 

//////////--------------------------------------------------------------------------------------------------------------=
//  calculation of X Axis speed using and position calculate regarding X_direction key or colision

always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN)
	begin
		Xspeed	<= INITIAL_X_SPEED;
		topLeftX_FixedPoint	<= INITIAL_X * FIXED_POINT_MULTIPLIER;
	end
	else begin
	
	// X collisions

	if (topLeftX_FixedPoint <= INITIAL_X* FIXED_POINT_MULTIPLIER) begin
		Xspeed <= INITIAL_X_SPEED;
	end
	if (topLeftX_FixedPoint >= x_FRAME_SIZE - 192* FIXED_POINT_MULTIPLIER) begin
		Xspeed <= -INITIAL_X_SPEED;
	end
	 
	
	if (startOfFrame == 1'b1 )
		topLeftX_FixedPoint  <= topLeftX_FixedPoint + Xspeed;
		//rope_speed	<= Xspeed;
					
	end
end

//get a better (64 times) resolution using integer   
assign 	topLeftX = topLeftX_FixedPoint / FIXED_POINT_MULTIPLIER ;   // note it must be 2^n 
assign 	topLeftY = topLeftY_FixedPoint / FIXED_POINT_MULTIPLIER ;    


endmodule
