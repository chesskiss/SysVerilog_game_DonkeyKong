// (c) Technion IIT, Department of Electrical Engineering 2021 
//-- Alex Grinshpun Apr 2017
//-- Dudy Nov 13 2017
// SystemVerilog version Alex Grinshpun May 2018
// coding convention dudy December 2018
// updaed Eyal Lev Feb 2021


module	monkey_moveCollision	(	
 
					input	logic	clk,
					input	logic	resetN,
					input	logic	startOfFrame,  // short pulse every start of frame 30Hz 
					input	logic	Y_up, 
					input	logic	Y_down,
					input	logic	X_right, 	
					input	logic	X_left,
					input logic collision_f_floor,
					input logic collision_f_ropes,// active in case of collision between two objects
					input logic collision_f_fruits,
					input logic collision_f_target,
					input logic collision_f_enemy,
					input logic collision_f_rope,
					input logic SingleHit_floor,
					input logic SingleHit_ropes,
					input logic SingleHit_fruits,
					input logic SingleHit_target,
					input logic SingleHit_enemy,
					input logic [3:0] HitEdgeCode,
					input logic [10:0] ropePixelX,
					input logic [10:0] ropePixelY,

					output	 logic signed 	[10:0]	topLeftX, // output the top left corner 
					output	 logic signed	[10:0]	topLeftY  // can be negative , if the object is partliy outside 
					
);


// a module used to generate the  ball trajectory.  

parameter int INITIAL_X = 32;
parameter int INITIAL_Y = 400;//128
parameter int INITIAL_X_SPEED = 0;
parameter int INITIAL_Y_SPEED = 0;
parameter int MAX_Y_SPEED = 230;
parameter int MAX_SPEED_X = 230;
const int  Y_ACCEL = -8;
const int  X_ACCEL = 200;
const int  Y_MOVE = 250;
const int  Y_MOVE_DOWN = 200;
const int  X_MOVE = 100; //


const int	FIXED_POINT_MULTIPLIER	=	64;
// FIXED_POINT_MULTIPLIER is used to enable working with integers in high resolution so that 
// we do all calculations with topLeftX_FixedPoint to get a resolution of 1/64 pixel in calcuatuions,
// we devide at the end by FIXED_POINT_MULTIPLIER which must be 2^n, to return to the initial proportions
const int	x_FRAME_SIZE	=	575 * FIXED_POINT_MULTIPLIER; // note it must be 2^n //639 ?
const int	y_FRAME_SIZE	=	479 * FIXED_POINT_MULTIPLIER;
const int	bracketOffset =	30;
const int   OBJECT_WIDTH_X = 64;

int Xspeed, topLeftX_FixedPoint; // local parameters 
int Yspeed, topLeftY_FixedPoint;

//////////--------------------------------------------------------------------------------------------------------------=
//  calculation 0f Y Axis speed using gravity or colision

always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin 
		Yspeed	<= INITIAL_Y_SPEED;
		topLeftY_FixedPoint	<= INITIAL_Y * FIXED_POINT_MULTIPLIER;
	end 
	else begin
	// colision Calcultaion 
		
			
		//hit bit map has one bit per edge:  Left-Top-Right-Bottom	 

		if(SingleHit_floor) begin
			if (HitEdgeCode [2] == 1 && Yspeed < 0)  // hit top border of brick  
					Yspeed <= -Yspeed; 	
			
				else if (HitEdgeCode [0] == 1 && Yspeed > 0 && Y_down != 1)// || (collision && HitEdgeCode [1] == 1 ))   hit bottom border of brick  
					Yspeed <= 0;
		end
				
				//else if ((HitEdgeCode [3] == 1 || HitEdgeCode [1] == 1))
					//Yspeed <= Yspeed;  //not redundent !
		
		// bottom collision
		if (topLeftY_FixedPoint > INITIAL_Y * FIXED_POINT_MULTIPLIER) begin
			topLeftY_FixedPoint <= INITIAL_Y * FIXED_POINT_MULTIPLIER;
			Yspeed <= 0;
		end
		
		// perform  position and speed integral only 30 times per second 
		
		if (startOfFrame == 1'b1) begin 
		
			topLeftY_FixedPoint  <= topLeftY_FixedPoint + Yspeed; // position interpolation 
				
			 // deAccelerate : slow the speed down every clock tick  
			if(topLeftY_FixedPoint < INITIAL_Y * FIXED_POINT_MULTIPLIER) begin
				if(collision_f_ropes == 1'b0 && collision_f_rope == 1'b0) begin
					if(Yspeed == Y_ACCEL)
						Yspeed <= Yspeed  - Y_ACCEL - 1 ;
					else
						Yspeed <= Yspeed  - Y_ACCEL ;
				end
				else
					Yspeed <= (Y_down && !Yspeed) ? (Yspeed + Y_MOVE_DOWN) : 0;
			
			end
			
			if (Y_up && !Yspeed) 
					Yspeed <= Yspeed - Y_MOVE  ;

			if (Y_down && !Yspeed && (topLeftY_FixedPoint > INITIAL_Y*FIXED_POINT_MULTIPLIER))
					Yspeed <= Yspeed + Y_MOVE  ;
					
			if (collision_f_enemy ||collision_f_target) begin
				topLeftY_FixedPoint	<= INITIAL_Y * FIXED_POINT_MULTIPLIER;
				// heart --;
			end
			
		end
	end
end 

//////////--------------------------------------------------------------------------------------------------------------=
//  calculation of X Axis speed using and position calculate regarding X_direction key or colision

always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN)
	begin
		Xspeed	<= INITIAL_X_SPEED;
		topLeftX_FixedPoint	<= INITIAL_X * FIXED_POINT_MULTIPLIER;
	end
	else begin

	
	// X collisions
	
	if (topLeftX_FixedPoint < 0) begin
		topLeftX_FixedPoint <= 0;
		Xspeed <= 0;
	end
	if (topLeftX_FixedPoint > x_FRAME_SIZE) begin
		topLeftX_FixedPoint <= x_FRAME_SIZE;
		Xspeed <= 0;
	end
	
	
	if (collision_f_rope && !X_left && !X_right && !ropePixelX[10] && (HitEdgeCode[3] || HitEdgeCode[2] || HitEdgeCode[1]))
					Xspeed <= 20;//ropePixelX;
	else if(collision_f_rope && !X_left && !X_right && ropePixelX[10] && (HitEdgeCode[3] || HitEdgeCode[2] || HitEdgeCode[1]))
					Xspeed <= -20;//-ropePixelX;
	
	
	if (startOfFrame == 1'b1 ) begin
	
	topLeftX_FixedPoint  <= topLeftX_FixedPoint + Xspeed;

	// X speed and deacceleration 
	
	if(Xspeed > 0) begin
		if(Xspeed < X_ACCEL)
			Xspeed <= 0;
		else
			Xspeed <= Xspeed  - X_ACCEL ;	
	end
	if(Xspeed < 0) begin
		if(Xspeed > -X_ACCEL)
			Xspeed <= 0;
		else
			Xspeed <= Xspeed  + X_ACCEL ;	
	end
	
	if (X_right && Xspeed < MAX_SPEED_X)  
				Xspeed <= Xspeed + X_MOVE; 

	if (X_left && Xspeed > (-MAX_SPEED_X))  
				Xspeed <= Xspeed - X_MOVE; 
					
	if (collision_f_enemy || collision_f_target)
					topLeftX_FixedPoint	<= INITIAL_X * FIXED_POINT_MULTIPLIER;	
	
		end // else begin
	end //ff begin
end

//get a better (64 times) resolution using integer   
assign 	topLeftX = topLeftX_FixedPoint / FIXED_POINT_MULTIPLIER ;   // note it must be 2^n 
assign 	topLeftY = topLeftY_FixedPoint / FIXED_POINT_MULTIPLIER ;    


endmodule
